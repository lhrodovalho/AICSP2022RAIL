* opamp voltage follower testbench

* Include SkyWater sky130 device models
.lib "/usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.param mc_mm_switch=0

.include "array.spice"
.include "ampa.spice"
.include "ampb.spice"
.include "params.spice"

VDD vdd 0 dc {pVDD}
VSS vss 0 0
ECM cm vss vdd vss 0.5

vin in cm dc 0 ac 1 PULSE({-pAMP} {pAMP} {pT/4} {pT*1m} {pT*1m} {pT/2} {pT})

iba vdd iba {pIB}
xa  oa in oa iba vdd vss ampa
ca  oa cm {pC}
ra  oa cm {pR}

ibb vdd ibb {pIB}
xb  ob in ob ibb vdd vss ampb
cb  ob cm {pC}
rb  ob cm {pR}

.option gmin=1e-15
*.option method=Gear
.tran {pT*1m} {pT}

.control

	run
	plot in oa ob
	wrdata ../data/ampa_vf_tran_step.txt in oa
	wrdata ../data/ampb_vf_tran_step.txt in ob
	
	let vmax = 2.5
	let vmin = 0.5
	let dv   = vmax-vmin
	
	meas tran slewpa trig v(oa) rise=1 val=vmin targ v(oa) rise=1 val=vmax
	meas tran slewma trig v(oa) fall=1 val=vmax targ v(oa) fall=1 val=vmin
	meas tran slewpb trig v(ob) rise=1 val=vmin targ v(ob) rise=1 val=vmax
	meas tran slewmb trig v(ob) fall=1 val=vmax targ v(ob) fall=1 val=vmin

	let slewrpa = dv/slewpa
	let slewrma = dv/slewma
	let slewrpb = dv/slewpb
	let slewrmb = dv/slewmb
	
	print slewrpa slewrma slewrpb slewrmb
	
.endc

.end
