* SPICE3 file created from pmos.ext - technology: sky130A

X0 a_2010_n960# a_1910_n990# a_1850_n960# w_n160_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=3e+11p pd=2.3e+06u as=3e+11p ps=2.3e+06u w=2e+06u l=500000u
X1 a_90_0# a_n10_n160# a_n80_0# w_n160_n80# sky130_fd_pr__pfet_g5v0d10v5 ad=3e+11p pd=2.3e+06u as=7e+11p ps=4.7e+06u w=2e+06u l=500000u
X2 a_730_n960# a_630_n990# a_570_n960# w_n160_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=3e+11p pd=2.3e+06u as=3e+11p ps=2.3e+06u w=2e+06u l=500000u
X3 a_890_n960# a_630_n990# a_730_n960# w_n160_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=3e+11p pd=2.3e+06u as=3e+11p ps=2.3e+06u w=2e+06u l=500000u
X4 a_2170_0# a_1910_n160# a_2010_0# w_n160_n80# sky130_fd_pr__pfet_g5v0d10v5 ad=3e+11p pd=2.3e+06u as=3e+11p ps=2.3e+06u w=2e+06u l=500000u
X5 a_90_n960# a_n10_n990# a_n80_n960# w_n160_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=3e+11p pd=2.3e+06u as=7e+11p ps=4.7e+06u w=2e+06u l=500000u
X6 a_1530_n960# a_1270_n990# a_1370_n960# w_n160_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=3e+11p pd=2.3e+06u as=3e+11p ps=2.3e+06u w=2e+06u l=500000u
X7 a_1690_n960# a_1590_n990# a_1530_n960# w_n160_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=3e+11p pd=2.3e+06u as=3e+11p ps=2.3e+06u w=2e+06u l=500000u
X8 a_1850_0# a_1590_n160# a_1690_0# w_n160_n80# sky130_fd_pr__pfet_g5v0d10v5 ad=3e+11p pd=2.3e+06u as=3e+11p ps=2.3e+06u w=2e+06u l=500000u
X9 a_2330_n960# a_2230_n990# a_2170_n960# w_n160_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=3e+11p pd=2.3e+06u as=3e+11p ps=2.3e+06u w=2e+06u l=500000u
X10 a_730_0# a_630_n160# a_570_0# w_n160_n80# sky130_fd_pr__pfet_g5v0d10v5 ad=3e+11p pd=2.3e+06u as=3e+11p ps=2.3e+06u w=2e+06u l=500000u
X11 a_2490_n960# a_2230_n990# a_2330_n960# w_n160_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=7e+11p pd=4.7e+06u as=3e+11p ps=2.3e+06u w=2e+06u l=500000u
X12 a_890_0# a_630_n160# a_730_0# w_n160_n80# sky130_fd_pr__pfet_g5v0d10v5 ad=3e+11p pd=2.3e+06u as=3e+11p ps=2.3e+06u w=2e+06u l=500000u
X13 a_250_n960# a_n10_n990# a_90_n960# w_n160_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=3e+11p pd=2.3e+06u as=3e+11p ps=2.3e+06u w=2e+06u l=500000u
X14 a_1210_0# a_950_n160# a_1050_0# w_n160_n80# sky130_fd_pr__pfet_g5v0d10v5 ad=3e+11p pd=2.3e+06u as=3e+11p ps=2.3e+06u w=2e+06u l=500000u
X15 a_1370_0# a_1270_n160# a_1210_0# w_n160_n80# sky130_fd_pr__pfet_g5v0d10v5 ad=3e+11p pd=2.3e+06u as=3e+11p ps=2.3e+06u w=2e+06u l=500000u
X16 a_250_0# a_n10_n160# a_90_0# w_n160_n80# sky130_fd_pr__pfet_g5v0d10v5 ad=3e+11p pd=2.3e+06u as=3e+11p ps=2.3e+06u w=2e+06u l=500000u
X17 a_2330_0# a_2230_n160# a_2170_0# w_n160_n80# sky130_fd_pr__pfet_g5v0d10v5 ad=3e+11p pd=2.3e+06u as=3e+11p ps=2.3e+06u w=2e+06u l=500000u
X18 a_1050_n960# a_950_n990# a_890_n960# w_n160_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=3e+11p pd=2.3e+06u as=3e+11p ps=2.3e+06u w=2e+06u l=500000u
X19 a_2490_0# a_2230_n160# a_2330_0# w_n160_n80# sky130_fd_pr__pfet_g5v0d10v5 ad=7e+11p pd=4.7e+06u as=3e+11p ps=2.3e+06u w=2e+06u l=500000u
X20 a_2010_0# a_1910_n160# a_1850_0# w_n160_n80# sky130_fd_pr__pfet_g5v0d10v5 ad=3e+11p pd=2.3e+06u as=3e+11p ps=2.3e+06u w=2e+06u l=500000u
X21 a_1850_n960# a_1590_n990# a_1690_n960# w_n160_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=3e+11p pd=2.3e+06u as=3e+11p ps=2.3e+06u w=2e+06u l=500000u
X22 a_1050_0# a_950_n160# a_890_0# w_n160_n80# sky130_fd_pr__pfet_g5v0d10v5 ad=3e+11p pd=2.3e+06u as=3e+11p ps=2.3e+06u w=2e+06u l=500000u
X23 a_410_n960# a_310_n990# a_250_n960# w_n160_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=3e+11p pd=2.3e+06u as=3e+11p ps=2.3e+06u w=2e+06u l=500000u
X24 a_570_n960# a_310_n990# a_410_n960# w_n160_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=3e+11p pd=2.3e+06u as=3e+11p ps=2.3e+06u w=2e+06u l=500000u
X25 a_410_0# a_310_n160# a_250_0# w_n160_n80# sky130_fd_pr__pfet_g5v0d10v5 ad=3e+11p pd=2.3e+06u as=3e+11p ps=2.3e+06u w=2e+06u l=500000u
X26 a_1530_0# a_1270_n160# a_1370_0# w_n160_n80# sky130_fd_pr__pfet_g5v0d10v5 ad=3e+11p pd=2.3e+06u as=3e+11p ps=2.3e+06u w=2e+06u l=500000u
X27 a_1210_n960# a_950_n990# a_1050_n960# w_n160_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=3e+11p pd=2.3e+06u as=3e+11p ps=2.3e+06u w=2e+06u l=500000u
X28 a_1370_n960# a_1270_n990# a_1210_n960# w_n160_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=3e+11p pd=2.3e+06u as=3e+11p ps=2.3e+06u w=2e+06u l=500000u
X29 a_2170_n960# a_1910_n990# a_2010_n960# w_n160_n1200# sky130_fd_pr__pfet_g5v0d10v5 ad=3e+11p pd=2.3e+06u as=3e+11p ps=2.3e+06u w=2e+06u l=500000u
X30 a_570_0# a_310_n160# a_410_0# w_n160_n80# sky130_fd_pr__pfet_g5v0d10v5 ad=3e+11p pd=2.3e+06u as=3e+11p ps=2.3e+06u w=2e+06u l=500000u
X31 a_1690_0# a_1590_n160# a_1530_0# w_n160_n80# sky130_fd_pr__pfet_g5v0d10v5 ad=3e+11p pd=2.3e+06u as=3e+11p ps=2.3e+06u w=2e+06u l=500000u
C0 w_n160_n1200# a_n80_n1360# 6.05fF **FLOATING
C1 w_n160_n80# a_n80_n1360# 6.05fF **FLOATING
