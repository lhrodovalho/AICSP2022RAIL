magic
tech sky130A
timestamp 1653815306
<< nwell >>
rect -80 -40 1320 320
rect -80 -600 1320 -240
<< mvpmos >>
rect -5 0 45 200
rect 75 0 125 200
rect 155 0 205 200
rect 235 0 285 200
rect 315 0 365 200
rect 395 0 445 200
rect 475 0 525 200
rect 555 0 605 200
rect 635 0 685 200
rect 715 0 765 200
rect 795 0 845 200
rect 875 0 925 200
rect 955 0 1005 200
rect 1035 0 1085 200
rect 1115 0 1165 200
rect 1195 0 1245 200
rect -5 -480 45 -280
rect 75 -480 125 -280
rect 155 -480 205 -280
rect 235 -480 285 -280
rect 315 -480 365 -280
rect 395 -480 445 -280
rect 475 -480 525 -280
rect 555 -480 605 -280
rect 635 -480 685 -280
rect 715 -480 765 -280
rect 795 -480 845 -280
rect 875 -480 925 -280
rect 955 -480 1005 -280
rect 1035 -480 1085 -280
rect 1115 -480 1165 -280
rect 1195 -480 1245 -280
<< mvpdiff >>
rect -40 189 -5 200
rect -40 171 -29 189
rect -11 171 -5 189
rect -40 149 -5 171
rect -40 131 -29 149
rect -11 131 -5 149
rect -40 109 -5 131
rect -40 91 -29 109
rect -11 91 -5 109
rect -40 69 -5 91
rect -40 51 -29 69
rect -11 51 -5 69
rect -40 29 -5 51
rect -40 11 -29 29
rect -11 11 -5 29
rect -40 0 -5 11
rect 45 189 75 200
rect 45 171 51 189
rect 69 171 75 189
rect 45 149 75 171
rect 45 131 51 149
rect 69 131 75 149
rect 45 109 75 131
rect 45 91 51 109
rect 69 91 75 109
rect 45 69 75 91
rect 45 51 51 69
rect 69 51 75 69
rect 45 29 75 51
rect 45 11 51 29
rect 69 11 75 29
rect 45 0 75 11
rect 125 189 155 200
rect 125 171 131 189
rect 149 171 155 189
rect 125 149 155 171
rect 125 131 131 149
rect 149 131 155 149
rect 125 109 155 131
rect 125 91 131 109
rect 149 91 155 109
rect 125 69 155 91
rect 125 51 131 69
rect 149 51 155 69
rect 125 29 155 51
rect 125 11 131 29
rect 149 11 155 29
rect 125 0 155 11
rect 205 189 235 200
rect 205 171 211 189
rect 229 171 235 189
rect 205 149 235 171
rect 205 131 211 149
rect 229 131 235 149
rect 205 109 235 131
rect 205 91 211 109
rect 229 91 235 109
rect 205 69 235 91
rect 205 51 211 69
rect 229 51 235 69
rect 205 29 235 51
rect 205 11 211 29
rect 229 11 235 29
rect 205 0 235 11
rect 285 189 315 200
rect 285 171 291 189
rect 309 171 315 189
rect 285 149 315 171
rect 285 131 291 149
rect 309 131 315 149
rect 285 109 315 131
rect 285 91 291 109
rect 309 91 315 109
rect 285 69 315 91
rect 285 51 291 69
rect 309 51 315 69
rect 285 29 315 51
rect 285 11 291 29
rect 309 11 315 29
rect 285 0 315 11
rect 365 189 395 200
rect 365 171 371 189
rect 389 171 395 189
rect 365 149 395 171
rect 365 131 371 149
rect 389 131 395 149
rect 365 109 395 131
rect 365 91 371 109
rect 389 91 395 109
rect 365 69 395 91
rect 365 51 371 69
rect 389 51 395 69
rect 365 29 395 51
rect 365 11 371 29
rect 389 11 395 29
rect 365 0 395 11
rect 445 189 475 200
rect 445 171 451 189
rect 469 171 475 189
rect 445 149 475 171
rect 445 131 451 149
rect 469 131 475 149
rect 445 109 475 131
rect 445 91 451 109
rect 469 91 475 109
rect 445 69 475 91
rect 445 51 451 69
rect 469 51 475 69
rect 445 29 475 51
rect 445 11 451 29
rect 469 11 475 29
rect 445 0 475 11
rect 525 189 555 200
rect 525 171 531 189
rect 549 171 555 189
rect 525 149 555 171
rect 525 131 531 149
rect 549 131 555 149
rect 525 109 555 131
rect 525 91 531 109
rect 549 91 555 109
rect 525 69 555 91
rect 525 51 531 69
rect 549 51 555 69
rect 525 29 555 51
rect 525 11 531 29
rect 549 11 555 29
rect 525 0 555 11
rect 605 189 635 200
rect 605 171 611 189
rect 629 171 635 189
rect 605 149 635 171
rect 605 131 611 149
rect 629 131 635 149
rect 605 109 635 131
rect 605 91 611 109
rect 629 91 635 109
rect 605 69 635 91
rect 605 51 611 69
rect 629 51 635 69
rect 605 29 635 51
rect 605 11 611 29
rect 629 11 635 29
rect 605 0 635 11
rect 685 189 715 200
rect 685 171 691 189
rect 709 171 715 189
rect 685 149 715 171
rect 685 131 691 149
rect 709 131 715 149
rect 685 109 715 131
rect 685 91 691 109
rect 709 91 715 109
rect 685 69 715 91
rect 685 51 691 69
rect 709 51 715 69
rect 685 29 715 51
rect 685 11 691 29
rect 709 11 715 29
rect 685 0 715 11
rect 765 189 795 200
rect 765 171 771 189
rect 789 171 795 189
rect 765 149 795 171
rect 765 131 771 149
rect 789 131 795 149
rect 765 109 795 131
rect 765 91 771 109
rect 789 91 795 109
rect 765 69 795 91
rect 765 51 771 69
rect 789 51 795 69
rect 765 29 795 51
rect 765 11 771 29
rect 789 11 795 29
rect 765 0 795 11
rect 845 189 875 200
rect 845 171 851 189
rect 869 171 875 189
rect 845 149 875 171
rect 845 131 851 149
rect 869 131 875 149
rect 845 109 875 131
rect 845 91 851 109
rect 869 91 875 109
rect 845 69 875 91
rect 845 51 851 69
rect 869 51 875 69
rect 845 29 875 51
rect 845 11 851 29
rect 869 11 875 29
rect 845 0 875 11
rect 925 189 955 200
rect 925 171 931 189
rect 949 171 955 189
rect 925 149 955 171
rect 925 131 931 149
rect 949 131 955 149
rect 925 109 955 131
rect 925 91 931 109
rect 949 91 955 109
rect 925 69 955 91
rect 925 51 931 69
rect 949 51 955 69
rect 925 29 955 51
rect 925 11 931 29
rect 949 11 955 29
rect 925 0 955 11
rect 1005 189 1035 200
rect 1005 171 1011 189
rect 1029 171 1035 189
rect 1005 149 1035 171
rect 1005 131 1011 149
rect 1029 131 1035 149
rect 1005 109 1035 131
rect 1005 91 1011 109
rect 1029 91 1035 109
rect 1005 69 1035 91
rect 1005 51 1011 69
rect 1029 51 1035 69
rect 1005 29 1035 51
rect 1005 11 1011 29
rect 1029 11 1035 29
rect 1005 0 1035 11
rect 1085 189 1115 200
rect 1085 171 1091 189
rect 1109 171 1115 189
rect 1085 149 1115 171
rect 1085 131 1091 149
rect 1109 131 1115 149
rect 1085 109 1115 131
rect 1085 91 1091 109
rect 1109 91 1115 109
rect 1085 69 1115 91
rect 1085 51 1091 69
rect 1109 51 1115 69
rect 1085 29 1115 51
rect 1085 11 1091 29
rect 1109 11 1115 29
rect 1085 0 1115 11
rect 1165 189 1195 200
rect 1165 171 1171 189
rect 1189 171 1195 189
rect 1165 149 1195 171
rect 1165 131 1171 149
rect 1189 131 1195 149
rect 1165 109 1195 131
rect 1165 91 1171 109
rect 1189 91 1195 109
rect 1165 69 1195 91
rect 1165 51 1171 69
rect 1189 51 1195 69
rect 1165 29 1195 51
rect 1165 11 1171 29
rect 1189 11 1195 29
rect 1165 0 1195 11
rect 1245 189 1280 200
rect 1245 171 1251 189
rect 1269 171 1280 189
rect 1245 149 1280 171
rect 1245 131 1251 149
rect 1269 131 1280 149
rect 1245 109 1280 131
rect 1245 91 1251 109
rect 1269 91 1280 109
rect 1245 69 1280 91
rect 1245 51 1251 69
rect 1269 51 1280 69
rect 1245 29 1280 51
rect 1245 11 1251 29
rect 1269 11 1280 29
rect 1245 0 1280 11
rect -40 -291 -5 -280
rect -40 -309 -29 -291
rect -11 -309 -5 -291
rect -40 -331 -5 -309
rect -40 -349 -29 -331
rect -11 -349 -5 -331
rect -40 -371 -5 -349
rect -40 -389 -29 -371
rect -11 -389 -5 -371
rect -40 -411 -5 -389
rect -40 -429 -29 -411
rect -11 -429 -5 -411
rect -40 -451 -5 -429
rect -40 -469 -29 -451
rect -11 -469 -5 -451
rect -40 -480 -5 -469
rect 45 -291 75 -280
rect 45 -309 51 -291
rect 69 -309 75 -291
rect 45 -331 75 -309
rect 45 -349 51 -331
rect 69 -349 75 -331
rect 45 -371 75 -349
rect 45 -389 51 -371
rect 69 -389 75 -371
rect 45 -411 75 -389
rect 45 -429 51 -411
rect 69 -429 75 -411
rect 45 -451 75 -429
rect 45 -469 51 -451
rect 69 -469 75 -451
rect 45 -480 75 -469
rect 125 -291 155 -280
rect 125 -309 131 -291
rect 149 -309 155 -291
rect 125 -331 155 -309
rect 125 -349 131 -331
rect 149 -349 155 -331
rect 125 -371 155 -349
rect 125 -389 131 -371
rect 149 -389 155 -371
rect 125 -411 155 -389
rect 125 -429 131 -411
rect 149 -429 155 -411
rect 125 -451 155 -429
rect 125 -469 131 -451
rect 149 -469 155 -451
rect 125 -480 155 -469
rect 205 -291 235 -280
rect 205 -309 211 -291
rect 229 -309 235 -291
rect 205 -331 235 -309
rect 205 -349 211 -331
rect 229 -349 235 -331
rect 205 -371 235 -349
rect 205 -389 211 -371
rect 229 -389 235 -371
rect 205 -411 235 -389
rect 205 -429 211 -411
rect 229 -429 235 -411
rect 205 -451 235 -429
rect 205 -469 211 -451
rect 229 -469 235 -451
rect 205 -480 235 -469
rect 285 -291 315 -280
rect 285 -309 291 -291
rect 309 -309 315 -291
rect 285 -331 315 -309
rect 285 -349 291 -331
rect 309 -349 315 -331
rect 285 -371 315 -349
rect 285 -389 291 -371
rect 309 -389 315 -371
rect 285 -411 315 -389
rect 285 -429 291 -411
rect 309 -429 315 -411
rect 285 -451 315 -429
rect 285 -469 291 -451
rect 309 -469 315 -451
rect 285 -480 315 -469
rect 365 -291 395 -280
rect 365 -309 371 -291
rect 389 -309 395 -291
rect 365 -331 395 -309
rect 365 -349 371 -331
rect 389 -349 395 -331
rect 365 -371 395 -349
rect 365 -389 371 -371
rect 389 -389 395 -371
rect 365 -411 395 -389
rect 365 -429 371 -411
rect 389 -429 395 -411
rect 365 -451 395 -429
rect 365 -469 371 -451
rect 389 -469 395 -451
rect 365 -480 395 -469
rect 445 -291 475 -280
rect 445 -309 451 -291
rect 469 -309 475 -291
rect 445 -331 475 -309
rect 445 -349 451 -331
rect 469 -349 475 -331
rect 445 -371 475 -349
rect 445 -389 451 -371
rect 469 -389 475 -371
rect 445 -411 475 -389
rect 445 -429 451 -411
rect 469 -429 475 -411
rect 445 -451 475 -429
rect 445 -469 451 -451
rect 469 -469 475 -451
rect 445 -480 475 -469
rect 525 -291 555 -280
rect 525 -309 531 -291
rect 549 -309 555 -291
rect 525 -331 555 -309
rect 525 -349 531 -331
rect 549 -349 555 -331
rect 525 -371 555 -349
rect 525 -389 531 -371
rect 549 -389 555 -371
rect 525 -411 555 -389
rect 525 -429 531 -411
rect 549 -429 555 -411
rect 525 -451 555 -429
rect 525 -469 531 -451
rect 549 -469 555 -451
rect 525 -480 555 -469
rect 605 -291 635 -280
rect 605 -309 611 -291
rect 629 -309 635 -291
rect 605 -331 635 -309
rect 605 -349 611 -331
rect 629 -349 635 -331
rect 605 -371 635 -349
rect 605 -389 611 -371
rect 629 -389 635 -371
rect 605 -411 635 -389
rect 605 -429 611 -411
rect 629 -429 635 -411
rect 605 -451 635 -429
rect 605 -469 611 -451
rect 629 -469 635 -451
rect 605 -480 635 -469
rect 685 -291 715 -280
rect 685 -309 691 -291
rect 709 -309 715 -291
rect 685 -331 715 -309
rect 685 -349 691 -331
rect 709 -349 715 -331
rect 685 -371 715 -349
rect 685 -389 691 -371
rect 709 -389 715 -371
rect 685 -411 715 -389
rect 685 -429 691 -411
rect 709 -429 715 -411
rect 685 -451 715 -429
rect 685 -469 691 -451
rect 709 -469 715 -451
rect 685 -480 715 -469
rect 765 -291 795 -280
rect 765 -309 771 -291
rect 789 -309 795 -291
rect 765 -331 795 -309
rect 765 -349 771 -331
rect 789 -349 795 -331
rect 765 -371 795 -349
rect 765 -389 771 -371
rect 789 -389 795 -371
rect 765 -411 795 -389
rect 765 -429 771 -411
rect 789 -429 795 -411
rect 765 -451 795 -429
rect 765 -469 771 -451
rect 789 -469 795 -451
rect 765 -480 795 -469
rect 845 -291 875 -280
rect 845 -309 851 -291
rect 869 -309 875 -291
rect 845 -331 875 -309
rect 845 -349 851 -331
rect 869 -349 875 -331
rect 845 -371 875 -349
rect 845 -389 851 -371
rect 869 -389 875 -371
rect 845 -411 875 -389
rect 845 -429 851 -411
rect 869 -429 875 -411
rect 845 -451 875 -429
rect 845 -469 851 -451
rect 869 -469 875 -451
rect 845 -480 875 -469
rect 925 -291 955 -280
rect 925 -309 931 -291
rect 949 -309 955 -291
rect 925 -331 955 -309
rect 925 -349 931 -331
rect 949 -349 955 -331
rect 925 -371 955 -349
rect 925 -389 931 -371
rect 949 -389 955 -371
rect 925 -411 955 -389
rect 925 -429 931 -411
rect 949 -429 955 -411
rect 925 -451 955 -429
rect 925 -469 931 -451
rect 949 -469 955 -451
rect 925 -480 955 -469
rect 1005 -291 1035 -280
rect 1005 -309 1011 -291
rect 1029 -309 1035 -291
rect 1005 -331 1035 -309
rect 1005 -349 1011 -331
rect 1029 -349 1035 -331
rect 1005 -371 1035 -349
rect 1005 -389 1011 -371
rect 1029 -389 1035 -371
rect 1005 -411 1035 -389
rect 1005 -429 1011 -411
rect 1029 -429 1035 -411
rect 1005 -451 1035 -429
rect 1005 -469 1011 -451
rect 1029 -469 1035 -451
rect 1005 -480 1035 -469
rect 1085 -291 1115 -280
rect 1085 -309 1091 -291
rect 1109 -309 1115 -291
rect 1085 -331 1115 -309
rect 1085 -349 1091 -331
rect 1109 -349 1115 -331
rect 1085 -371 1115 -349
rect 1085 -389 1091 -371
rect 1109 -389 1115 -371
rect 1085 -411 1115 -389
rect 1085 -429 1091 -411
rect 1109 -429 1115 -411
rect 1085 -451 1115 -429
rect 1085 -469 1091 -451
rect 1109 -469 1115 -451
rect 1085 -480 1115 -469
rect 1165 -291 1195 -280
rect 1165 -309 1171 -291
rect 1189 -309 1195 -291
rect 1165 -331 1195 -309
rect 1165 -349 1171 -331
rect 1189 -349 1195 -331
rect 1165 -371 1195 -349
rect 1165 -389 1171 -371
rect 1189 -389 1195 -371
rect 1165 -411 1195 -389
rect 1165 -429 1171 -411
rect 1189 -429 1195 -411
rect 1165 -451 1195 -429
rect 1165 -469 1171 -451
rect 1189 -469 1195 -451
rect 1165 -480 1195 -469
rect 1245 -291 1280 -280
rect 1245 -309 1251 -291
rect 1269 -309 1280 -291
rect 1245 -331 1280 -309
rect 1245 -349 1251 -331
rect 1269 -349 1280 -331
rect 1245 -371 1280 -349
rect 1245 -389 1251 -371
rect 1269 -389 1280 -371
rect 1245 -411 1280 -389
rect 1245 -429 1251 -411
rect 1269 -429 1280 -411
rect 1245 -451 1280 -429
rect 1245 -469 1251 -451
rect 1269 -469 1280 -451
rect 1245 -480 1280 -469
<< mvpdiffc >>
rect -29 171 -11 189
rect -29 131 -11 149
rect -29 91 -11 109
rect -29 51 -11 69
rect -29 11 -11 29
rect 51 171 69 189
rect 51 131 69 149
rect 51 91 69 109
rect 51 51 69 69
rect 51 11 69 29
rect 131 171 149 189
rect 131 131 149 149
rect 131 91 149 109
rect 131 51 149 69
rect 131 11 149 29
rect 211 171 229 189
rect 211 131 229 149
rect 211 91 229 109
rect 211 51 229 69
rect 211 11 229 29
rect 291 171 309 189
rect 291 131 309 149
rect 291 91 309 109
rect 291 51 309 69
rect 291 11 309 29
rect 371 171 389 189
rect 371 131 389 149
rect 371 91 389 109
rect 371 51 389 69
rect 371 11 389 29
rect 451 171 469 189
rect 451 131 469 149
rect 451 91 469 109
rect 451 51 469 69
rect 451 11 469 29
rect 531 171 549 189
rect 531 131 549 149
rect 531 91 549 109
rect 531 51 549 69
rect 531 11 549 29
rect 611 171 629 189
rect 611 131 629 149
rect 611 91 629 109
rect 611 51 629 69
rect 611 11 629 29
rect 691 171 709 189
rect 691 131 709 149
rect 691 91 709 109
rect 691 51 709 69
rect 691 11 709 29
rect 771 171 789 189
rect 771 131 789 149
rect 771 91 789 109
rect 771 51 789 69
rect 771 11 789 29
rect 851 171 869 189
rect 851 131 869 149
rect 851 91 869 109
rect 851 51 869 69
rect 851 11 869 29
rect 931 171 949 189
rect 931 131 949 149
rect 931 91 949 109
rect 931 51 949 69
rect 931 11 949 29
rect 1011 171 1029 189
rect 1011 131 1029 149
rect 1011 91 1029 109
rect 1011 51 1029 69
rect 1011 11 1029 29
rect 1091 171 1109 189
rect 1091 131 1109 149
rect 1091 91 1109 109
rect 1091 51 1109 69
rect 1091 11 1109 29
rect 1171 171 1189 189
rect 1171 131 1189 149
rect 1171 91 1189 109
rect 1171 51 1189 69
rect 1171 11 1189 29
rect 1251 171 1269 189
rect 1251 131 1269 149
rect 1251 91 1269 109
rect 1251 51 1269 69
rect 1251 11 1269 29
rect -29 -309 -11 -291
rect -29 -349 -11 -331
rect -29 -389 -11 -371
rect -29 -429 -11 -411
rect -29 -469 -11 -451
rect 51 -309 69 -291
rect 51 -349 69 -331
rect 51 -389 69 -371
rect 51 -429 69 -411
rect 51 -469 69 -451
rect 131 -309 149 -291
rect 131 -349 149 -331
rect 131 -389 149 -371
rect 131 -429 149 -411
rect 131 -469 149 -451
rect 211 -309 229 -291
rect 211 -349 229 -331
rect 211 -389 229 -371
rect 211 -429 229 -411
rect 211 -469 229 -451
rect 291 -309 309 -291
rect 291 -349 309 -331
rect 291 -389 309 -371
rect 291 -429 309 -411
rect 291 -469 309 -451
rect 371 -309 389 -291
rect 371 -349 389 -331
rect 371 -389 389 -371
rect 371 -429 389 -411
rect 371 -469 389 -451
rect 451 -309 469 -291
rect 451 -349 469 -331
rect 451 -389 469 -371
rect 451 -429 469 -411
rect 451 -469 469 -451
rect 531 -309 549 -291
rect 531 -349 549 -331
rect 531 -389 549 -371
rect 531 -429 549 -411
rect 531 -469 549 -451
rect 611 -309 629 -291
rect 611 -349 629 -331
rect 611 -389 629 -371
rect 611 -429 629 -411
rect 611 -469 629 -451
rect 691 -309 709 -291
rect 691 -349 709 -331
rect 691 -389 709 -371
rect 691 -429 709 -411
rect 691 -469 709 -451
rect 771 -309 789 -291
rect 771 -349 789 -331
rect 771 -389 789 -371
rect 771 -429 789 -411
rect 771 -469 789 -451
rect 851 -309 869 -291
rect 851 -349 869 -331
rect 851 -389 869 -371
rect 851 -429 869 -411
rect 851 -469 869 -451
rect 931 -309 949 -291
rect 931 -349 949 -331
rect 931 -389 949 -371
rect 931 -429 949 -411
rect 931 -469 949 -451
rect 1011 -309 1029 -291
rect 1011 -349 1029 -331
rect 1011 -389 1029 -371
rect 1011 -429 1029 -411
rect 1011 -469 1029 -451
rect 1091 -309 1109 -291
rect 1091 -349 1109 -331
rect 1091 -389 1109 -371
rect 1091 -429 1109 -411
rect 1091 -469 1109 -451
rect 1171 -309 1189 -291
rect 1171 -349 1189 -331
rect 1171 -389 1189 -371
rect 1171 -429 1189 -411
rect 1171 -469 1189 -451
rect 1251 -309 1269 -291
rect 1251 -349 1269 -331
rect 1251 -389 1269 -371
rect 1251 -429 1269 -411
rect 1251 -469 1269 -451
<< mvpsubdiff >>
rect -40 360 1280 400
rect -40 -680 1280 -640
<< mvnsubdiff >>
rect -40 240 1280 280
rect -40 -560 1280 -520
<< poly >>
rect -5 200 45 215
rect 75 200 125 215
rect 155 200 205 215
rect 235 200 285 215
rect 315 200 365 215
rect 395 200 445 215
rect 475 200 525 215
rect 555 200 605 215
rect 635 200 685 215
rect 715 200 765 215
rect 795 200 845 215
rect 875 200 925 215
rect 955 200 1005 215
rect 1035 200 1085 215
rect 1115 200 1165 215
rect 1195 200 1245 215
rect -5 -40 45 0
rect 75 -40 125 0
rect -5 -80 125 -40
rect 155 -40 205 0
rect 235 -40 285 0
rect 155 -80 285 -40
rect 315 -40 365 0
rect 395 -40 445 0
rect 315 -80 445 -40
rect 475 -40 525 0
rect 555 -40 605 0
rect 475 -80 605 -40
rect 635 -40 685 0
rect 715 -40 765 0
rect 635 -80 765 -40
rect 795 -40 845 0
rect 875 -40 925 0
rect 795 -80 925 -40
rect 955 -40 1005 0
rect 1035 -40 1085 0
rect 955 -80 1085 -40
rect 1115 -40 1165 0
rect 1195 -40 1245 0
rect 1115 -80 1245 -40
rect -5 -240 125 -200
rect -5 -280 45 -240
rect 75 -280 125 -240
rect 155 -240 285 -200
rect 155 -280 205 -240
rect 235 -280 285 -240
rect 315 -240 445 -200
rect 315 -280 365 -240
rect 395 -280 445 -240
rect 475 -240 605 -200
rect 475 -280 525 -240
rect 555 -280 605 -240
rect 635 -240 765 -200
rect 635 -280 685 -240
rect 715 -280 765 -240
rect 795 -240 925 -200
rect 795 -280 845 -240
rect 875 -280 925 -240
rect 955 -240 1085 -200
rect 955 -280 1005 -240
rect 1035 -280 1085 -240
rect 1115 -240 1245 -200
rect 1115 -280 1165 -240
rect 1195 -280 1245 -240
rect -5 -495 45 -480
rect 75 -495 125 -480
rect 155 -495 205 -480
rect 235 -495 285 -480
rect 315 -495 365 -480
rect 395 -495 445 -480
rect 475 -495 525 -480
rect 555 -495 605 -480
rect 635 -495 685 -480
rect 715 -495 765 -480
rect 795 -495 845 -480
rect 875 -495 925 -480
rect 955 -495 1005 -480
rect 1035 -495 1085 -480
rect 1115 -495 1165 -480
rect 1195 -495 1245 -480
<< locali >>
rect -40 189 0 200
rect -40 171 -29 189
rect -11 171 0 189
rect -40 149 0 171
rect -40 131 -29 149
rect -11 131 0 149
rect -40 109 0 131
rect -40 91 -29 109
rect -11 91 0 109
rect -40 69 0 91
rect -40 51 -29 69
rect -11 51 0 69
rect -40 29 0 51
rect -40 11 -29 29
rect -11 11 0 29
rect -40 0 0 11
rect 40 189 80 200
rect 40 171 51 189
rect 69 171 80 189
rect 40 149 80 171
rect 40 131 51 149
rect 69 131 80 149
rect 40 109 80 131
rect 40 91 51 109
rect 69 91 80 109
rect 40 69 80 91
rect 40 51 51 69
rect 69 51 80 69
rect 40 29 80 51
rect 40 11 51 29
rect 69 11 80 29
rect 40 0 80 11
rect 120 189 160 200
rect 120 171 131 189
rect 149 171 160 189
rect 120 149 160 171
rect 120 131 131 149
rect 149 131 160 149
rect 120 109 160 131
rect 120 91 131 109
rect 149 91 160 109
rect 120 69 160 91
rect 120 51 131 69
rect 149 51 160 69
rect 120 29 160 51
rect 120 11 131 29
rect 149 11 160 29
rect 120 0 160 11
rect 200 189 240 200
rect 200 171 211 189
rect 229 171 240 189
rect 200 149 240 171
rect 200 131 211 149
rect 229 131 240 149
rect 200 109 240 131
rect 200 91 211 109
rect 229 91 240 109
rect 200 69 240 91
rect 200 51 211 69
rect 229 51 240 69
rect 200 29 240 51
rect 200 11 211 29
rect 229 11 240 29
rect 200 0 240 11
rect 280 189 320 200
rect 280 171 291 189
rect 309 171 320 189
rect 280 149 320 171
rect 280 131 291 149
rect 309 131 320 149
rect 280 109 320 131
rect 280 91 291 109
rect 309 91 320 109
rect 280 69 320 91
rect 280 51 291 69
rect 309 51 320 69
rect 280 29 320 51
rect 280 11 291 29
rect 309 11 320 29
rect 280 0 320 11
rect 360 189 400 200
rect 360 171 371 189
rect 389 171 400 189
rect 360 149 400 171
rect 360 131 371 149
rect 389 131 400 149
rect 360 109 400 131
rect 360 91 371 109
rect 389 91 400 109
rect 360 69 400 91
rect 360 51 371 69
rect 389 51 400 69
rect 360 29 400 51
rect 360 11 371 29
rect 389 11 400 29
rect 360 0 400 11
rect 440 189 480 200
rect 440 171 451 189
rect 469 171 480 189
rect 440 149 480 171
rect 440 131 451 149
rect 469 131 480 149
rect 440 109 480 131
rect 440 91 451 109
rect 469 91 480 109
rect 440 69 480 91
rect 440 51 451 69
rect 469 51 480 69
rect 440 29 480 51
rect 440 11 451 29
rect 469 11 480 29
rect 440 0 480 11
rect 520 189 560 200
rect 520 171 531 189
rect 549 171 560 189
rect 520 149 560 171
rect 520 131 531 149
rect 549 131 560 149
rect 520 109 560 131
rect 520 91 531 109
rect 549 91 560 109
rect 520 69 560 91
rect 520 51 531 69
rect 549 51 560 69
rect 520 29 560 51
rect 520 11 531 29
rect 549 11 560 29
rect 520 0 560 11
rect 600 189 640 200
rect 600 171 611 189
rect 629 171 640 189
rect 600 149 640 171
rect 600 131 611 149
rect 629 131 640 149
rect 600 109 640 131
rect 600 91 611 109
rect 629 91 640 109
rect 600 69 640 91
rect 600 51 611 69
rect 629 51 640 69
rect 600 29 640 51
rect 600 11 611 29
rect 629 11 640 29
rect 600 0 640 11
rect 680 189 720 200
rect 680 171 691 189
rect 709 171 720 189
rect 680 149 720 171
rect 680 131 691 149
rect 709 131 720 149
rect 680 109 720 131
rect 680 91 691 109
rect 709 91 720 109
rect 680 69 720 91
rect 680 51 691 69
rect 709 51 720 69
rect 680 29 720 51
rect 680 11 691 29
rect 709 11 720 29
rect 680 0 720 11
rect 760 189 800 200
rect 760 171 771 189
rect 789 171 800 189
rect 760 149 800 171
rect 760 131 771 149
rect 789 131 800 149
rect 760 109 800 131
rect 760 91 771 109
rect 789 91 800 109
rect 760 69 800 91
rect 760 51 771 69
rect 789 51 800 69
rect 760 29 800 51
rect 760 11 771 29
rect 789 11 800 29
rect 760 0 800 11
rect 840 189 880 200
rect 840 171 851 189
rect 869 171 880 189
rect 840 149 880 171
rect 840 131 851 149
rect 869 131 880 149
rect 840 109 880 131
rect 840 91 851 109
rect 869 91 880 109
rect 840 69 880 91
rect 840 51 851 69
rect 869 51 880 69
rect 840 29 880 51
rect 840 11 851 29
rect 869 11 880 29
rect 840 0 880 11
rect 920 189 960 200
rect 920 171 931 189
rect 949 171 960 189
rect 920 149 960 171
rect 920 131 931 149
rect 949 131 960 149
rect 920 109 960 131
rect 920 91 931 109
rect 949 91 960 109
rect 920 69 960 91
rect 920 51 931 69
rect 949 51 960 69
rect 920 29 960 51
rect 920 11 931 29
rect 949 11 960 29
rect 920 0 960 11
rect 1000 189 1040 200
rect 1000 171 1011 189
rect 1029 171 1040 189
rect 1000 149 1040 171
rect 1000 131 1011 149
rect 1029 131 1040 149
rect 1000 109 1040 131
rect 1000 91 1011 109
rect 1029 91 1040 109
rect 1000 69 1040 91
rect 1000 51 1011 69
rect 1029 51 1040 69
rect 1000 29 1040 51
rect 1000 11 1011 29
rect 1029 11 1040 29
rect 1000 0 1040 11
rect 1080 189 1120 200
rect 1080 171 1091 189
rect 1109 171 1120 189
rect 1080 149 1120 171
rect 1080 131 1091 149
rect 1109 131 1120 149
rect 1080 109 1120 131
rect 1080 91 1091 109
rect 1109 91 1120 109
rect 1080 69 1120 91
rect 1080 51 1091 69
rect 1109 51 1120 69
rect 1080 29 1120 51
rect 1080 11 1091 29
rect 1109 11 1120 29
rect 1080 0 1120 11
rect 1160 189 1200 200
rect 1160 171 1171 189
rect 1189 171 1200 189
rect 1160 149 1200 171
rect 1160 131 1171 149
rect 1189 131 1200 149
rect 1160 109 1200 131
rect 1160 91 1171 109
rect 1189 91 1200 109
rect 1160 69 1200 91
rect 1160 51 1171 69
rect 1189 51 1200 69
rect 1160 29 1200 51
rect 1160 11 1171 29
rect 1189 11 1200 29
rect 1160 0 1200 11
rect 1240 189 1280 200
rect 1240 171 1251 189
rect 1269 171 1280 189
rect 1240 149 1280 171
rect 1240 131 1251 149
rect 1269 131 1280 149
rect 1240 109 1280 131
rect 1240 91 1251 109
rect 1269 91 1280 109
rect 1240 69 1280 91
rect 1240 51 1251 69
rect 1269 51 1280 69
rect 1240 29 1280 51
rect 1240 11 1251 29
rect 1269 11 1280 29
rect 1240 0 1280 11
rect 0 -80 280 -40
rect 320 -80 600 -40
rect 640 -80 920 -40
rect 960 -80 1240 -40
rect 0 -240 280 -200
rect 320 -240 600 -200
rect 640 -240 920 -200
rect 960 -240 1240 -200
rect -40 -291 0 -280
rect -40 -309 -29 -291
rect -11 -309 0 -291
rect -40 -331 0 -309
rect -40 -349 -29 -331
rect -11 -349 0 -331
rect -40 -371 0 -349
rect -40 -389 -29 -371
rect -11 -389 0 -371
rect -40 -411 0 -389
rect -40 -429 -29 -411
rect -11 -429 0 -411
rect -40 -451 0 -429
rect -40 -469 -29 -451
rect -11 -469 0 -451
rect -40 -480 0 -469
rect 40 -291 80 -280
rect 40 -309 51 -291
rect 69 -309 80 -291
rect 40 -331 80 -309
rect 40 -349 51 -331
rect 69 -349 80 -331
rect 40 -371 80 -349
rect 40 -389 51 -371
rect 69 -389 80 -371
rect 40 -411 80 -389
rect 40 -429 51 -411
rect 69 -429 80 -411
rect 40 -451 80 -429
rect 40 -469 51 -451
rect 69 -469 80 -451
rect 40 -480 80 -469
rect 120 -291 160 -280
rect 120 -309 131 -291
rect 149 -309 160 -291
rect 120 -331 160 -309
rect 120 -349 131 -331
rect 149 -349 160 -331
rect 120 -371 160 -349
rect 120 -389 131 -371
rect 149 -389 160 -371
rect 120 -411 160 -389
rect 120 -429 131 -411
rect 149 -429 160 -411
rect 120 -451 160 -429
rect 120 -469 131 -451
rect 149 -469 160 -451
rect 120 -480 160 -469
rect 200 -291 240 -280
rect 200 -309 211 -291
rect 229 -309 240 -291
rect 200 -331 240 -309
rect 200 -349 211 -331
rect 229 -349 240 -331
rect 200 -371 240 -349
rect 200 -389 211 -371
rect 229 -389 240 -371
rect 200 -411 240 -389
rect 200 -429 211 -411
rect 229 -429 240 -411
rect 200 -451 240 -429
rect 200 -469 211 -451
rect 229 -469 240 -451
rect 200 -480 240 -469
rect 280 -291 320 -280
rect 280 -309 291 -291
rect 309 -309 320 -291
rect 280 -331 320 -309
rect 280 -349 291 -331
rect 309 -349 320 -331
rect 280 -371 320 -349
rect 280 -389 291 -371
rect 309 -389 320 -371
rect 280 -411 320 -389
rect 280 -429 291 -411
rect 309 -429 320 -411
rect 280 -451 320 -429
rect 280 -469 291 -451
rect 309 -469 320 -451
rect 280 -480 320 -469
rect 360 -291 400 -280
rect 360 -309 371 -291
rect 389 -309 400 -291
rect 360 -331 400 -309
rect 360 -349 371 -331
rect 389 -349 400 -331
rect 360 -371 400 -349
rect 360 -389 371 -371
rect 389 -389 400 -371
rect 360 -411 400 -389
rect 360 -429 371 -411
rect 389 -429 400 -411
rect 360 -451 400 -429
rect 360 -469 371 -451
rect 389 -469 400 -451
rect 360 -480 400 -469
rect 440 -291 480 -280
rect 440 -309 451 -291
rect 469 -309 480 -291
rect 440 -331 480 -309
rect 440 -349 451 -331
rect 469 -349 480 -331
rect 440 -371 480 -349
rect 440 -389 451 -371
rect 469 -389 480 -371
rect 440 -411 480 -389
rect 440 -429 451 -411
rect 469 -429 480 -411
rect 440 -451 480 -429
rect 440 -469 451 -451
rect 469 -469 480 -451
rect 440 -480 480 -469
rect 520 -291 560 -280
rect 520 -309 531 -291
rect 549 -309 560 -291
rect 520 -331 560 -309
rect 520 -349 531 -331
rect 549 -349 560 -331
rect 520 -371 560 -349
rect 520 -389 531 -371
rect 549 -389 560 -371
rect 520 -411 560 -389
rect 520 -429 531 -411
rect 549 -429 560 -411
rect 520 -451 560 -429
rect 520 -469 531 -451
rect 549 -469 560 -451
rect 520 -480 560 -469
rect 600 -291 640 -280
rect 600 -309 611 -291
rect 629 -309 640 -291
rect 600 -331 640 -309
rect 600 -349 611 -331
rect 629 -349 640 -331
rect 600 -371 640 -349
rect 600 -389 611 -371
rect 629 -389 640 -371
rect 600 -411 640 -389
rect 600 -429 611 -411
rect 629 -429 640 -411
rect 600 -451 640 -429
rect 600 -469 611 -451
rect 629 -469 640 -451
rect 600 -480 640 -469
rect 680 -291 720 -280
rect 680 -309 691 -291
rect 709 -309 720 -291
rect 680 -331 720 -309
rect 680 -349 691 -331
rect 709 -349 720 -331
rect 680 -371 720 -349
rect 680 -389 691 -371
rect 709 -389 720 -371
rect 680 -411 720 -389
rect 680 -429 691 -411
rect 709 -429 720 -411
rect 680 -451 720 -429
rect 680 -469 691 -451
rect 709 -469 720 -451
rect 680 -480 720 -469
rect 760 -291 800 -280
rect 760 -309 771 -291
rect 789 -309 800 -291
rect 760 -331 800 -309
rect 760 -349 771 -331
rect 789 -349 800 -331
rect 760 -371 800 -349
rect 760 -389 771 -371
rect 789 -389 800 -371
rect 760 -411 800 -389
rect 760 -429 771 -411
rect 789 -429 800 -411
rect 760 -451 800 -429
rect 760 -469 771 -451
rect 789 -469 800 -451
rect 760 -480 800 -469
rect 840 -291 880 -280
rect 840 -309 851 -291
rect 869 -309 880 -291
rect 840 -331 880 -309
rect 840 -349 851 -331
rect 869 -349 880 -331
rect 840 -371 880 -349
rect 840 -389 851 -371
rect 869 -389 880 -371
rect 840 -411 880 -389
rect 840 -429 851 -411
rect 869 -429 880 -411
rect 840 -451 880 -429
rect 840 -469 851 -451
rect 869 -469 880 -451
rect 840 -480 880 -469
rect 920 -291 960 -280
rect 920 -309 931 -291
rect 949 -309 960 -291
rect 920 -331 960 -309
rect 920 -349 931 -331
rect 949 -349 960 -331
rect 920 -371 960 -349
rect 920 -389 931 -371
rect 949 -389 960 -371
rect 920 -411 960 -389
rect 920 -429 931 -411
rect 949 -429 960 -411
rect 920 -451 960 -429
rect 920 -469 931 -451
rect 949 -469 960 -451
rect 920 -480 960 -469
rect 1000 -291 1040 -280
rect 1000 -309 1011 -291
rect 1029 -309 1040 -291
rect 1000 -331 1040 -309
rect 1000 -349 1011 -331
rect 1029 -349 1040 -331
rect 1000 -371 1040 -349
rect 1000 -389 1011 -371
rect 1029 -389 1040 -371
rect 1000 -411 1040 -389
rect 1000 -429 1011 -411
rect 1029 -429 1040 -411
rect 1000 -451 1040 -429
rect 1000 -469 1011 -451
rect 1029 -469 1040 -451
rect 1000 -480 1040 -469
rect 1080 -291 1120 -280
rect 1080 -309 1091 -291
rect 1109 -309 1120 -291
rect 1080 -331 1120 -309
rect 1080 -349 1091 -331
rect 1109 -349 1120 -331
rect 1080 -371 1120 -349
rect 1080 -389 1091 -371
rect 1109 -389 1120 -371
rect 1080 -411 1120 -389
rect 1080 -429 1091 -411
rect 1109 -429 1120 -411
rect 1080 -451 1120 -429
rect 1080 -469 1091 -451
rect 1109 -469 1120 -451
rect 1080 -480 1120 -469
rect 1160 -291 1200 -280
rect 1160 -309 1171 -291
rect 1189 -309 1200 -291
rect 1160 -331 1200 -309
rect 1160 -349 1171 -331
rect 1189 -349 1200 -331
rect 1160 -371 1200 -349
rect 1160 -389 1171 -371
rect 1189 -389 1200 -371
rect 1160 -411 1200 -389
rect 1160 -429 1171 -411
rect 1189 -429 1200 -411
rect 1160 -451 1200 -429
rect 1160 -469 1171 -451
rect 1189 -469 1200 -451
rect 1160 -480 1200 -469
rect 1240 -291 1280 -280
rect 1240 -309 1251 -291
rect 1269 -309 1280 -291
rect 1240 -331 1280 -309
rect 1240 -349 1251 -331
rect 1269 -349 1280 -331
rect 1240 -371 1280 -349
rect 1240 -389 1251 -371
rect 1269 -389 1280 -371
rect 1240 -411 1280 -389
rect 1240 -429 1251 -411
rect 1269 -429 1280 -411
rect 1240 -451 1280 -429
rect 1240 -469 1251 -451
rect 1269 -469 1280 -451
rect 1240 -480 1280 -469
<< metal1 >>
rect -40 -80 0 200
rect 120 -80 160 -40
rect 280 -80 320 40
rect 440 -80 480 40
rect 600 -80 640 200
rect 760 -80 800 -40
rect 920 -80 960 40
rect 1080 -80 1120 40
rect 1240 -80 1280 200
rect -40 -480 0 -200
rect 120 -240 160 -200
rect 280 -320 320 -200
rect 440 -320 480 -200
rect 600 -480 640 -200
rect 760 -240 800 -200
rect 920 -320 960 -200
rect 1080 -320 1120 -200
rect 1240 -480 1280 -200
<< metal2 >>
rect -40 160 1280 200
rect 40 0 560 40
rect 680 0 1200 40
rect -80 -160 1320 -120
rect 40 -320 560 -280
rect 680 -320 1200 -280
rect -40 -480 1280 -440
<< end >>
