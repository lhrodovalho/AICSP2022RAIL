magic
tech sky130A
timestamp 1653735127
<< nwell >>
rect -120 -200 720 320
<< mvpmos >>
rect -5 0 45 200
rect 75 0 125 200
rect 155 0 205 200
rect 235 0 285 200
rect 315 0 365 200
rect 395 0 445 200
rect 475 0 525 200
rect 555 0 605 200
<< mvpdiff >>
rect -40 189 -5 200
rect -40 171 -29 189
rect -11 171 -5 189
rect -40 149 -5 171
rect -40 131 -29 149
rect -11 131 -5 149
rect -40 109 -5 131
rect -40 91 -29 109
rect -11 91 -5 109
rect -40 0 -5 91
rect 45 109 75 200
rect 45 91 51 109
rect 69 91 75 109
rect 45 69 75 91
rect 45 51 51 69
rect 69 51 75 69
rect 45 29 75 51
rect 45 11 51 29
rect 69 11 75 29
rect 45 0 75 11
rect 125 189 155 200
rect 125 171 131 189
rect 149 171 155 189
rect 125 149 155 171
rect 125 131 131 149
rect 149 131 155 149
rect 125 109 155 131
rect 125 91 131 109
rect 149 91 155 109
rect 125 0 155 91
rect 205 109 235 200
rect 205 91 211 109
rect 229 91 235 109
rect 205 69 235 91
rect 205 51 211 69
rect 229 51 235 69
rect 205 29 235 51
rect 205 11 211 29
rect 229 11 235 29
rect 205 0 235 11
rect 285 189 315 200
rect 285 171 291 189
rect 309 171 315 189
rect 285 149 315 171
rect 285 131 291 149
rect 309 131 315 149
rect 285 109 315 131
rect 285 91 291 109
rect 309 91 315 109
rect 285 0 315 91
rect 365 109 395 200
rect 365 91 371 109
rect 389 91 395 109
rect 365 69 395 91
rect 365 51 371 69
rect 389 51 395 69
rect 365 29 395 51
rect 365 11 371 29
rect 389 11 395 29
rect 365 0 395 11
rect 445 189 475 200
rect 445 171 451 189
rect 469 171 475 189
rect 445 149 475 171
rect 445 131 451 149
rect 469 131 475 149
rect 445 109 475 131
rect 445 91 451 109
rect 469 91 475 109
rect 445 0 475 91
rect 525 109 555 200
rect 525 91 531 109
rect 549 91 555 109
rect 525 69 555 91
rect 525 51 531 69
rect 549 51 555 69
rect 525 29 555 51
rect 525 11 531 29
rect 549 11 555 29
rect 525 0 555 11
rect 605 189 640 200
rect 605 171 611 189
rect 629 171 640 189
rect 605 149 640 171
rect 605 131 611 149
rect 629 131 640 149
rect 605 109 640 131
rect 605 91 611 109
rect 629 91 640 109
rect 605 0 640 91
<< mvpdiffc >>
rect -29 171 -11 189
rect -29 131 -11 149
rect -29 91 -11 109
rect 51 91 69 109
rect 51 51 69 69
rect 51 11 69 29
rect 131 171 149 189
rect 131 131 149 149
rect 131 91 149 109
rect 211 91 229 109
rect 211 51 229 69
rect 211 11 229 29
rect 291 171 309 189
rect 291 131 309 149
rect 291 91 309 109
rect 371 91 389 109
rect 371 51 389 69
rect 371 11 389 29
rect 451 171 469 189
rect 451 131 469 149
rect 451 91 469 109
rect 531 91 549 109
rect 531 51 549 69
rect 531 11 549 29
rect 611 171 629 189
rect 611 131 629 149
rect 611 91 629 109
<< mvpsubdiff >>
rect -80 360 680 400
rect -80 -280 680 -240
<< mvnsubdiff >>
rect -80 240 680 280
rect -80 -160 680 -120
<< poly >>
rect -5 200 45 215
rect 75 200 125 215
rect 155 200 205 215
rect 235 200 285 215
rect 315 200 365 215
rect 395 200 445 215
rect 475 200 525 215
rect 555 200 605 215
rect -5 -40 45 0
rect 75 -40 125 0
rect -5 -80 125 -40
rect 155 -40 205 0
rect 235 -40 285 0
rect 155 -80 285 -40
rect 315 -40 365 0
rect 395 -40 445 0
rect 315 -80 445 -40
rect 475 -40 525 0
rect 555 -40 605 0
rect 475 -80 605 -40
<< locali >>
rect -40 189 640 200
rect -40 171 -29 189
rect -11 171 131 189
rect 149 171 291 189
rect 309 171 451 189
rect 469 171 611 189
rect 629 171 640 189
rect -40 160 640 171
rect -40 149 0 160
rect -40 131 -29 149
rect -11 131 0 149
rect -40 109 0 131
rect 120 149 160 160
rect 120 131 131 149
rect 149 131 160 149
rect -40 91 -29 109
rect -11 91 0 109
rect -40 80 0 91
rect 40 109 80 120
rect 40 91 51 109
rect 69 91 80 109
rect 40 69 80 91
rect 120 109 160 131
rect 280 149 320 160
rect 280 131 291 149
rect 309 131 320 149
rect 120 91 131 109
rect 149 91 160 109
rect 120 80 160 91
rect 200 109 240 120
rect 200 91 211 109
rect 229 91 240 109
rect 40 51 51 69
rect 69 51 80 69
rect 40 40 80 51
rect 200 69 240 91
rect 280 109 320 131
rect 440 149 480 160
rect 440 131 451 149
rect 469 131 480 149
rect 280 91 291 109
rect 309 91 320 109
rect 280 80 320 91
rect 360 109 400 120
rect 360 91 371 109
rect 389 91 400 109
rect 200 51 211 69
rect 229 51 240 69
rect 200 40 240 51
rect 360 69 400 91
rect 440 109 480 131
rect 600 149 640 160
rect 600 131 611 149
rect 629 131 640 149
rect 440 91 451 109
rect 469 91 480 109
rect 440 80 480 91
rect 520 109 560 120
rect 520 91 531 109
rect 549 91 560 109
rect 360 51 371 69
rect 389 51 400 69
rect 360 40 400 51
rect 520 69 560 91
rect 600 109 640 131
rect 600 91 611 109
rect 629 91 640 109
rect 600 80 640 91
rect 520 51 531 69
rect 549 51 560 69
rect 520 40 560 51
rect 40 29 560 40
rect 40 11 51 29
rect 69 11 211 29
rect 229 11 371 29
rect 389 11 531 29
rect 549 11 560 29
rect 40 0 560 11
rect 40 -80 560 -40
<< end >>
